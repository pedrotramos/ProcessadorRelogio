
LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY memoriaROM IS
    GENERIC (
        dataWidth : NATURAL := 18;
        addrWidth : NATURAL := 10
    );
    PORT (
        Endereco : IN std_logic_vector (addrWidth - 1 DOWNTO 0);
        Dado     : OUT std_logic_vector (dataWidth - 1 DOWNTO 0)
    );
END ENTITY;

ARCHITECTURE assincrona OF memoriaROM IS

    TYPE blocoMemoria IS ARRAY(0 TO 2 ** addrWidth - 1) OF std_logic_vector(dataWidth - 1 DOWNTO 0);

    FUNCTION initMemory
        RETURN blocoMemoria IS VARIABLE tmp : blocoMemoria := (OTHERS => (OTHERS => '0'));
    BEGIN
        tmp(0)   := b"111101010000000000";
        tmp(1)   := b"111101100000000000";
        tmp(2)   := b"111101110000000000";
        tmp(3)   := b"111110000000000000";
        tmp(4)   := b"111110010000000000";
        tmp(5)   := b"111000000000000000";
        tmp(6)   := b"111000000000000000";
        tmp(7)   := b"111000010000000000";
        tmp(8)   := b"111000100000000000";
        tmp(9)   := b"111000110000000000";
        tmp(10)  := b"111001000000000000";
        tmp(11)  := b"111001010000000000";
        tmp(12)  := b"111001100000000010";
        tmp(13)  := b"111001110000000001";
        tmp(14)  := b"111010000000001100";
        tmp(15)  := b"111010010000001010";
        tmp(16)  := b"100100010000000010";
        tmp(17)  := b"000100010000000001";
        tmp(18)  := b"110000000001100111";
        tmp(19)  := b"100100100000000001";
        tmp(20)  := b"000100100000000001";
        tmp(21)  := b"110000000010101000";
        tmp(22)  := b"100100000000000000";
        tmp(23)  := b"000100000000000000";
        tmp(24)  := b"110000000000011011";
        tmp(25)  := b"000100000000000001";
        tmp(26)  := b"110000000000100010";
        tmp(27)  := b"101000000000001110";
        tmp(28)  := b"101000010000001111";
        tmp(29)  := b"101000100000010000";
        tmp(30)  := b"101000110000010001";
        tmp(31)  := b"101001000000010010";
        tmp(32)  := b"101001010000010011";
        tmp(33)  := b"001000000011011101";
        tmp(34)  := b"101010010000001110";
        tmp(35)  := b"101010000000001111";
        tmp(36)  := b"101000100000010000";
        tmp(37)  := b"101000110000010001";
        tmp(38)  := b"101001000000010010";
        tmp(39)  := b"101001010000010011";
        tmp(40)  := b"001000000011011101";
        tmp(41)  := b"100101000000010100";
        tmp(42)  := b"000101000000000001";
        tmp(43)  := b"110000000000101101";
        tmp(44)  := b"001000000000010000";
        tmp(45)  := b"100101000000010101";
        tmp(46)  := b"000000000000001001";
        tmp(47)  := b"110000000000110010";
        tmp(48)  := b"010000000000000001";
        tmp(49)  := b"001000000000010000";
        tmp(50)  := b"111000000000000000";
        tmp(51)  := b"000000010000000101";
        tmp(52)  := b"110000000000110111";
        tmp(53)  := b"010000010000000001";
        tmp(54)  := b"001000000000010000";
        tmp(55)  := b"111000010000000000";
        tmp(56)  := b"000000100000001001";
        tmp(57)  := b"110000000000111100";
        tmp(58)  := b"010000100000000001";
        tmp(59)  := b"001000000000010000";
        tmp(60)  := b"111000100000000000";
        tmp(61)  := b"000000110000000101";
        tmp(62)  := b"110000000001000001";
        tmp(63)  := b"010000110000000001";
        tmp(64)  := b"001000000000010000";
        tmp(65)  := b"111000110000000000";
        tmp(66)  := b"000001100000000001";
        tmp(67)  := b"110000000001000111";
        tmp(68)  := b"000001100000000010";
        tmp(69)  := b"110000000001001011";
        tmp(70)  := b"001000000001011010";
        tmp(71)  := b"000001110000000001";
        tmp(72)  := b"110000000001001111";
        tmp(73)  := b"010001100000000001";
        tmp(74)  := b"001000000001100000";
        tmp(75)  := b"000001110000000001";
        tmp(76)  := b"110000000001010100";
        tmp(77)  := b"010001100000000001";
        tmp(78)  := b"001000000001100000";
        tmp(79)  := b"000010010000001111";
        tmp(80)  := b"110000000000000000";
        tmp(81)  := b"010001100000000001";
        tmp(82)  := b"111010010000001111";
        tmp(83)  := b"001000000001100000";
        tmp(84)  := b"000010010000001111";
        tmp(85)  := b"110000000000000000";
        tmp(86)  := b"111001100000000001";
        tmp(87)  := b"111001110000000000";
        tmp(88)  := b"111010010000001111";
        tmp(89)  := b"001000000001100000";
        tmp(90)  := b"000001100000001001";
        tmp(91)  := b"110000000001011110";
        tmp(92)  := b"010001100000000001";
        tmp(93)  := b"001000000001100000";
        tmp(94)  := b"111001100000000000";
        tmp(95)  := b"010001010000000001";
        tmp(96)  := b"000001000000001001";
        tmp(97)  := b"110000000001100100";
        tmp(98)  := b"010001000000000001";
        tmp(99)  := b"001000000000010000";
        tmp(100) := b"111001000000000000";
        tmp(101) := b"010001010000000001";
        tmp(102) := b"001000000000010000";
        tmp(103) := b"100000010000001010";
        tmp(104) := b"000000010000000000";
        tmp(105) := b"110000000010100010";
        tmp(106) := b"100000100000001011";
        tmp(107) := b"000000100000000000";
        tmp(108) := b"110000000010011100";
        tmp(109) := b"100000110000001100";
        tmp(110) := b"000000110000000000";
        tmp(111) := b"110000000010000101";
        tmp(112) := b"100001000000001101";
        tmp(113) := b"000001000000000000";
        tmp(114) := b"110000000001110100";
        tmp(115) := b"001000000000010110";
        tmp(116) := b"000001010000000010";
        tmp(117) := b"110000000001111011";
        tmp(118) := b"010001010000000001";
        tmp(119) := b"000001110000000001";
        tmp(120) := b"110000000001111101";
        tmp(121) := b"010001110000000001";
        tmp(122) := b"001000000000010110";
        tmp(123) := b"111001010000000000";
        tmp(124) := b"001000000001110111";
        tmp(125) := b"011001110000000001";
        tmp(126) := b"000010010000001111";
        tmp(127) := b"110000000010000001";
        tmp(128) := b"001000000010000011";
        tmp(129) := b"111010010000001010";
        tmp(130) := b"001000000000010110";
        tmp(131) := b"111010010000001111";
        tmp(132) := b"001000000000010110";
        tmp(133) := b"000001000000001001";
        tmp(134) := b"110000000010011000";
        tmp(135) := b"000001000000000011";
        tmp(136) := b"110000000010010000";
        tmp(137) := b"010001000000000001";
        tmp(138) := b"000001100000001001";
        tmp(139) := b"110000000010011010";
        tmp(140) := b"000001100000000010";
        tmp(141) := b"110000000010010100";
        tmp(142) := b"010001100000000001";
        tmp(143) := b"001000000000010110";
        tmp(144) := b"000001010000000010";
        tmp(145) := b"110000000010011000";
        tmp(146) := b"010001000000000001";
        tmp(147) := b"001000000010001010";
        tmp(148) := b"000001110000000001";
        tmp(149) := b"110000000010011000";
        tmp(150) := b"010001100000000001";
        tmp(151) := b"001000000000010110";
        tmp(152) := b"111001000000000000";
        tmp(153) := b"001000000010001010";
        tmp(154) := b"111001100000000001";
        tmp(155) := b"001000000000010110";
        tmp(156) := b"000000110000000101";
        tmp(157) := b"110000000010100000";
        tmp(158) := b"010000110000000001";
        tmp(159) := b"001000000000010110";
        tmp(160) := b"111000110000000000";
        tmp(161) := b"001000000000010110";
        tmp(162) := b"000000100000001001";
        tmp(163) := b"110000000010100110";
        tmp(164) := b"010000100000000001";
        tmp(165) := b"001000000000010110";
        tmp(166) := b"111000100000000000";
        tmp(167) := b"001000000000010110";
        tmp(168) := b"100000010000001010";
        tmp(169) := b"000000010000000000";
        tmp(170) := b"110000000010110101";
        tmp(171) := b"100000100000001011";
        tmp(172) := b"000000100000000000";
        tmp(173) := b"110000000011000000";
        tmp(174) := b"100000110000001100";
        tmp(175) := b"000000110000000000";
        tmp(176) := b"110000000011001011";
        tmp(177) := b"100001000000001101";
        tmp(178) := b"000001000000000000";
        tmp(179) := b"110000000011011101";
        tmp(180) := b"001000000011010110";
        tmp(181) := b"000101010000001001";
        tmp(182) := b"110000000010111001";
        tmp(183) := b"010101010000000001";
        tmp(184) := b"001000000011010110";
        tmp(185) := b"111101010000000000";
        tmp(186) := b"000101100000000101";
        tmp(187) := b"110000000010111110";
        tmp(188) := b"010101100000000001";
        tmp(189) := b"001000000011010110";
        tmp(190) := b"111101100000000000";
        tmp(191) := b"001000000011010110";
        tmp(192) := b"000101110000001001";
        tmp(193) := b"110000000011000100";
        tmp(194) := b"010101110000000001";
        tmp(195) := b"001000000011010110";
        tmp(196) := b"111101110000000000";
        tmp(197) := b"000110000000000101";
        tmp(198) := b"110000000011001001";
        tmp(199) := b"010110000000000001";
        tmp(200) := b"001000000011010110";
        tmp(201) := b"111110000000000000";
        tmp(202) := b"001000000011010110";
        tmp(203) := b"000110010000001001";
        tmp(204) := b"110000000011001111";
        tmp(205) := b"010110010000000001";
        tmp(206) := b"001000000011010110";
        tmp(207) := b"111110010000000000";
        tmp(208) := b"000000000000001001";
        tmp(209) := b"110000000011010100";
        tmp(210) := b"010000000000000001";
        tmp(211) := b"001000000011010110";
        tmp(212) := b"111000000000000000";
        tmp(213) := b"001000000011010110";
        tmp(214) := b"101101010000001110";
        tmp(215) := b"101101100000001111";
        tmp(216) := b"101101110000010000";
        tmp(217) := b"101110000000010001";
        tmp(218) := b"101110010000010010";
        tmp(219) := b"101000000000010011";
        tmp(220) := b"001000000011011101";
        tmp(221) := b"100101000000010100";
        tmp(222) := b"000101000000000001";
        tmp(223) := b"110000000011100001";
        tmp(224) := b"001000000000010000";
        tmp(225) := b"100101000000010101";
        tmp(226) := b"000101010000000000";
        tmp(227) := b"110000000011100110";
        tmp(228) := b"011101010000000001";
        tmp(229) := b"001000000000101101";
        tmp(230) := b"111101010000001001";
        tmp(231) := b"000101100000000000";
        tmp(232) := b"110000000011101011";
        tmp(233) := b"011101100000000001";
        tmp(234) := b"001000000000101101";
        tmp(235) := b"111101100000000101";
        tmp(236) := b"000101110000000000";
        tmp(237) := b"110000000011110000";
        tmp(238) := b"011101110000000001";
        tmp(239) := b"001000000000101101";
        tmp(240) := b"111101110000001001";
        tmp(241) := b"000110000000000000";
        tmp(242) := b"110000000011110101";
        tmp(243) := b"011110000000000001";
        tmp(244) := b"001000000000101101";
        tmp(245) := b"111110000000000101";
        tmp(246) := b"000110010000000000";
        tmp(247) := b"110000000011111010";
        tmp(248) := b"011110010000000001";
        tmp(249) := b"001000000000101101";
        tmp(250) := b"111110010000001001";
        tmp(251) := b"011000000000000001";
        tmp(252) := b"001000000000101101";

        RETURN tmp;
    END initMemory;

    SIGNAL memROM : blocoMemoria := initMemory;

BEGIN
    Dado <= memROM (to_integer(unsigned(Endereco)));
END ARCHITECTURE;