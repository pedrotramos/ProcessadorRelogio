
        LIBRARY IEEE;
        USE IEEE.std_logic_1164.ALL;
        USE ieee.numeric_std.ALL;

        ENTITY memoriaROM IS
            GENERIC (
                dataWidth : NATURAL := 17;
                addrWidth : NATURAL := 10
            );
            PORT (
                Endereco : IN std_logic_vector (addrWidth - 1 DOWNTO 0);
                Dado     : OUT std_logic_vector (dataWidth - 1 DOWNTO 0)
            );
        END ENTITY;

        ARCHITECTURE assincrona OF memoriaROM IS

            TYPE blocoMemoria IS ARRAY(0 TO 2 ** addrWidth - 1) OF std_logic_vector(dataWidth - 1 DOWNTO 0);

            FUNCTION initMemory
                RETURN blocoMemoria IS VARIABLE tmp : blocoMemoria := (OTHERS => (OTHERS => '0'));
            BEGIN
        tmp(0):= b"111011110000000000";
tmp(1):= b"111100000000000000";
tmp(2):= b"111100010000000000";
tmp(3):= b"111100100000000000";
tmp(4):= b"111100110000000000";
tmp(5):= b"111101000000000000";
tmp(6):= b"111000000000000000";
tmp(7):= b"111000010000000000";
tmp(8):= b"111000100000000000";
tmp(9):= b"111000110000000000";
tmp(10):= b"111001000000000000";
tmp(11):= b"111001010000000000";
tmp(12):= b"111001100000000010";
tmp(13):= b"111001110000000001";
tmp(14):= b"111010000000001100";
tmp(15):= b"111010010000001010";
tmp(16):= b"100110010000000100";
tmp(17):= b"000110010000000001";
tmp(18):= b"110000000100010010";
tmp(19):= b"100011000000000011";
tmp(20):= b"000011000000000001";
tmp(21):= b"110000000010111010";
tmp(22):= b"100010110000000010";
tmp(23):= b"000010110000000001";
tmp(24):= b"110000000001100111";
tmp(25):= b"100010100000000001";
tmp(26):= b"000010100000000000";
tmp(27):= b"110000000000011110";
tmp(28):= b"000010100000000001";
tmp(29):= b"110000000000100101";
tmp(30):= b"101000000000001110";
tmp(31):= b"101000010000001111";
tmp(32):= b"101000100000010000";
tmp(33):= b"101000110000010001";
tmp(34):= b"101001000000010010";
tmp(35):= b"101001010000010011";
tmp(36):= b"001000000000101100";
tmp(37):= b"101010010000001110";
tmp(38):= b"101010000000001111";
tmp(39):= b"101000100000010000";
tmp(40):= b"101000110000010001";
tmp(41):= b"101001100000010010";
tmp(42):= b"101001110000010011";
tmp(43):= b"001000000000101100";
tmp(44):= b"100011100000010100";
tmp(45):= b"000011100000000001";
tmp(46):= b"110000000000110000";
tmp(47):= b"001000000000010000";
tmp(48):= b"100011100000010101";
tmp(49):= b"000000000000001001";
tmp(50):= b"110000000000110101";
tmp(51):= b"010000000000000001";
tmp(52):= b"001000000000010000";
tmp(53):= b"111000000000000000";
tmp(54):= b"000000010000000101";
tmp(55):= b"110000000000111010";
tmp(56):= b"010000010000000001";
tmp(57):= b"001000000000010000";
tmp(58):= b"111000010000000000";
tmp(59):= b"000000100000001001";
tmp(60):= b"110000000000111111";
tmp(61):= b"010000100000000001";
tmp(62):= b"001000000000010000";
tmp(63):= b"111000100000000000";
tmp(64):= b"000000110000000101";
tmp(65):= b"110000000001000100";
tmp(66):= b"010000110000000001";
tmp(67):= b"001000000000010000";
tmp(68):= b"111000110000000000";
tmp(69):= b"000001100000000001";
tmp(70):= b"110000000001001010";
tmp(71):= b"000001100000000010";
tmp(72):= b"110000000001001110";
tmp(73):= b"001000000001011010";
tmp(74):= b"000001110000000001";
tmp(75):= b"110000000001010010";
tmp(76):= b"010001100000000001";
tmp(77):= b"001000000001100000";
tmp(78):= b"000001110000000001";
tmp(79):= b"110000000001010111";
tmp(80):= b"010001100000000001";
tmp(81):= b"001000000001100000";
tmp(82):= b"000010010000001111";
tmp(83):= b"110000000000000110";
tmp(84):= b"010001100000000001";
tmp(85):= b"111010010000001111";
tmp(86):= b"001000000001100000";
tmp(87):= b"111001100000000001";
tmp(88):= b"111001110000000000";
tmp(89):= b"001000000001100000";
tmp(90):= b"000001100000001001";
tmp(91):= b"110000000001011110";
tmp(92):= b"010001100000000001";
tmp(93):= b"001000000001100000";
tmp(94):= b"111001100000000000";
tmp(95):= b"010001110000000001";
tmp(96):= b"000001000000001001";
tmp(97):= b"110000000001100100";
tmp(98):= b"010001000000000001";
tmp(99):= b"001000000000010000";
tmp(100):= b"111001000000000000";
tmp(101):= b"010001010000000001";
tmp(102):= b"001000000000010000";
tmp(103):= b"100101010000001010";
tmp(104):= b"000101010000000000";
tmp(105):= b"110000000001110001";
tmp(106):= b"100101100000001011";
tmp(107):= b"000101100000000000";
tmp(108):= b"110000000001111000";
tmp(109):= b"100101110000001100";
tmp(110):= b"000101110000000000";
tmp(111):= b"110000000001111111";
tmp(112):= b"001000000000011001";
tmp(113):= b"100101010000001010";
tmp(114):= b"000101010000000001";
tmp(115):= b"110000000010000110";
tmp(116):= b"100011100000010100";
tmp(117):= b"000011100000000001";
tmp(118):= b"110000000010000110";
tmp(119):= b"001000000001110001";
tmp(120):= b"100101100000001011";
tmp(121):= b"000101100000000001";
tmp(122):= b"110000000010001100";
tmp(123):= b"100011100000010100";
tmp(124):= b"000011100000000001";
tmp(125):= b"110000000010001100";
tmp(126):= b"001000000001111000";
tmp(127):= b"100101110000001100";
tmp(128):= b"000101110000000001";
tmp(129):= b"110000000010010010";
tmp(130):= b"100011100000010100";
tmp(131):= b"000011100000000001";
tmp(132):= b"110000000010010010";
tmp(133):= b"001000000001111111";
tmp(134):= b"000000100000001001";
tmp(135):= b"110000000010001010";
tmp(136):= b"010000100000000001";
tmp(137):= b"001000000000011001";
tmp(138):= b"111000100000000000";
tmp(139):= b"001000000000011001";
tmp(140):= b"000000110000000101";
tmp(141):= b"110000000010010000";
tmp(142):= b"010000110000000001";
tmp(143):= b"001000000000011001";
tmp(144):= b"111000110000000000";
tmp(145):= b"001000000000011001";
tmp(146):= b"000001100000000001";
tmp(147):= b"110000000010010111";
tmp(148):= b"000001100000000010";
tmp(149):= b"110000000010011011";
tmp(150):= b"001000000010100111";
tmp(151):= b"000001110000000001";
tmp(152):= b"110000000010011111";
tmp(153):= b"010001100000000001";
tmp(154):= b"001000000010101101";
tmp(155):= b"000001110000000001";
tmp(156):= b"110000000010100100";
tmp(157):= b"010001100000000001";
tmp(158):= b"001000000010101101";
tmp(159):= b"000010010000001111";
tmp(160):= b"110000000010110100";
tmp(161):= b"010001100000000001";
tmp(162):= b"111010010000001111";
tmp(163):= b"001000000010101101";
tmp(164):= b"111001100000000001";
tmp(165):= b"111001110000000000";
tmp(166):= b"001000000010101101";
tmp(167):= b"000001100000001001";
tmp(168):= b"110000000010101011";
tmp(169):= b"010001100000000001";
tmp(170):= b"001000000010101101";
tmp(171):= b"111001100000000000";
tmp(172):= b"010001110000000001";
tmp(173):= b"000001000000001001";
tmp(174):= b"110000000010110001";
tmp(175):= b"010001000000000001";
tmp(176):= b"001000000000011001";
tmp(177):= b"111001000000000000";
tmp(178):= b"010001010000000001";
tmp(179):= b"001000000000011001";
tmp(180):= b"111001000000000000";
tmp(181):= b"111001010000000000";
tmp(182):= b"111001100000000010";
tmp(183):= b"111001110000000001";
tmp(184):= b"111010010000001010";
tmp(185):= b"001000000000011001";
tmp(186):= b"100101010000001010";
tmp(187):= b"000101010000000000";
tmp(188):= b"110000000011000111";
tmp(189):= b"100101100000001011";
tmp(190):= b"000101100000000000";
tmp(191):= b"110000000011001110";
tmp(192):= b"100101110000001100";
tmp(193):= b"000101110000000000";
tmp(194):= b"110000000011010101";
tmp(195):= b"100110000000001101";
tmp(196):= b"000110000000000000";
tmp(197):= b"110000000011011100";
tmp(198):= b"001000000100001011";
tmp(199):= b"100101010000001010";
tmp(200):= b"000101010000000001";
tmp(201):= b"110000000011100011";
tmp(202):= b"100011100000010100";
tmp(203):= b"000011100000000001";
tmp(204):= b"110000000011100011";
tmp(205):= b"001000000011000111";
tmp(206):= b"100101100000001011";
tmp(207):= b"000101100000000001";
tmp(208):= b"110000000011101110";
tmp(209):= b"100011100000010100";
tmp(210):= b"000011100000000001";
tmp(211):= b"110000000011101110";
tmp(212):= b"001000000011001110";
tmp(213):= b"100101110000001100";
tmp(214):= b"000101110000000001";
tmp(215):= b"110000000011111001";
tmp(216):= b"100011100000010100";
tmp(217):= b"000011100000000001";
tmp(218):= b"110000000011111001";
tmp(219):= b"001000000011010101";
tmp(220):= b"100110000000001101";
tmp(221):= b"000110000000000001";
tmp(222):= b"110000000100000100";
tmp(223):= b"100011100000010100";
tmp(224):= b"000011100000000001";
tmp(225):= b"110000000100000100";
tmp(226):= b"001000000011011100";
tmp(227):= b"000011110000001001";
tmp(228):= b"110000000011100111";
tmp(229):= b"010011110000000001";
tmp(230):= b"001000000100001011";
tmp(231):= b"111011110000000000";
tmp(232):= b"000100000000000101";
tmp(233):= b"110000000011101100";
tmp(234):= b"010100000000000001";
tmp(235):= b"001000000100001011";
tmp(236):= b"111100000000000000";
tmp(237):= b"001000000100001011";
tmp(238):= b"000100010000001001";
tmp(239):= b"110000000011110010";
tmp(240):= b"010100010000000001";
tmp(241):= b"001000000100001011";
tmp(242):= b"111100010000000000";
tmp(243):= b"000100100000000101";
tmp(244):= b"110000000011110111";
tmp(245):= b"010100100000000001";
tmp(246):= b"001000000100001011";
tmp(247):= b"111100100000000000";
tmp(248):= b"001000000100001011";
tmp(249):= b"000100110000001001";
tmp(250):= b"110000000011111101";
tmp(251):= b"010100110000000001";
tmp(252):= b"001000000100001011";
tmp(253):= b"111100110000000000";
tmp(254):= b"000101000000001001";
tmp(255):= b"110000000100000010";
tmp(256):= b"010101000000000001";
tmp(257):= b"001000000100001011";
tmp(258):= b"111101000000000000";
tmp(259):= b"001000000100001011";
tmp(260):= b"111011110000000000";
tmp(261):= b"111100000000000000";
tmp(262):= b"111100010000000000";
tmp(263):= b"111100100000000000";
tmp(264):= b"111100110000000000";
tmp(265):= b"111101000000000000";
tmp(266):= b"001000000100001011";
tmp(267):= b"101011110000001110";
tmp(268):= b"101100000000001111";
tmp(269):= b"101100010000010000";
tmp(270):= b"101100100000010001";
tmp(271):= b"101100110000010010";
tmp(272):= b"101101000000010011";
tmp(273):= b"001000000000101100";
tmp(274):= b"101011110000001110";
tmp(275):= b"101100000000001111";
tmp(276):= b"101100010000010000";
tmp(277):= b"101100100000010001";
tmp(278):= b"101100110000010010";
tmp(279):= b"101101000000010011";
tmp(280):= b"100011100000010100";
tmp(281):= b"000011100000000001";
tmp(282):= b"110000000100011100";
tmp(283):= b"001000000100011000";
tmp(284):= b"100011100000010101";
tmp(285):= b"000011110000000000";
tmp(286):= b"110000000100100001";
tmp(287):= b"011011110000000001";
tmp(288):= b"001000000101000001";
tmp(289):= b"111011110000001001";
tmp(290):= b"000100000000000000";
tmp(291):= b"110000000100100110";
tmp(292):= b"011100000000000001";
tmp(293):= b"001000000101000001";
tmp(294):= b"111100000000000101";
tmp(295):= b"000100010000000000";
tmp(296):= b"110000000100101011";
tmp(297):= b"011100010000000001";
tmp(298):= b"001000000101000001";
tmp(299):= b"111100010000001001";
tmp(300):= b"000100100000000000";
tmp(301):= b"110000000100110000";
tmp(302):= b"011100100000000001";
tmp(303):= b"001000000101000001";
tmp(304):= b"111100100000000101";
tmp(305):= b"000100110000000000";
tmp(306):= b"110000000100110101";
tmp(307):= b"011100110000000001";
tmp(308):= b"001000000101000001";
tmp(309):= b"000101000000000000";
tmp(310):= b"110000000100111010";
tmp(311):= b"111100110000001001";
tmp(312):= b"011101000000000001";
tmp(313):= b"001000000101000001";
tmp(314):= b"111011110000000000";
tmp(315):= b"111100000000000000";
tmp(316):= b"111100010000000000";
tmp(317):= b"111100100000000000";
tmp(318):= b"111100110000000000";
tmp(319):= b"111101000000000000";
tmp(320):= b"001000000101000001";
tmp(321):= b"101011110000001110";
tmp(322):= b"101100000000001111";
tmp(323):= b"101100010000010000";
tmp(324):= b"101100100000010001";
tmp(325):= b"101100110000010010";
tmp(326):= b"101101000000010011";
tmp(327):= b"001000000000110001";

            RETURN tmp;
        END initMemory;

        SIGNAL memROM : blocoMemoria := initMemory;

        BEGIN
            Dado <= memROM (to_integer(unsigned(Endereco)));
        END ARCHITECTURE;
        